module lab2(a, b, c, d, f1, f2, f3, f4, f5, f6, f7):
  input a, b, c, d;
  output f1, f2, f3, f4, f5, f6, f7;
  assign f1 = something;f
endmodule
