module question1(a, b, c);

    input a, b;
    output c;

    n

endmodule